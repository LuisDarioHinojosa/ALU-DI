`timescale 1ns / 1ps

module ALUA_TB;

	reg[7:0] A;
	reg[7:0] B;
	reg [1:0] S;
	wire [7:0]IS;
	wire cout;

	ALUA uut (
		.A(A), 
		.B(B), 
		.S(S), 
		.IS(IS),
		.cout(cout)
	);

	initial begin


	#100;
	A = 8'b00001111;
	B = 8'b00000101;
	S = 0;
	#100;

	#100;
	A = 8'b00001111;
	B = 8'b00000101;
	S = 1;
	#100;



	#100;
	A = 8'b00001111;
	B = 8'b00000101;
	S = 2;
	#100;

	#100;
	A = 8'b00001111;
	B = 8'b00000101;
	S = 3;
	#100;




/*
 	 // AND TB
	#100;
	A = 0;
	B = 0;
	S = 0;
	#100;


	#100;
	A = 0;
	B = 1;
	S = 0;
	#100;


	#100;
	A = 1;
	B = 0;
	S = 0;
	#100;


	#100;
	A = 1;
	B = 1;
	S = 0;
	#100;



	// OR TB 
	
	#100;
	A = 0;
	B = 0;
	S = 1;
	#100;


	#100;
	A = 0;
	B = 1;
	S = 1;
	#100;


	#100;
	A = 1;
	B = 0;
	S = 1;
	#100;


	#100;
	A = 1;
	B = 1;
	S = 1;
	#100;



	// XOR TB 
	
	#100;
	A = 0;
	B = 0;
	S = 2;
	#100;


	#100;
	A = 0;
	B = 1;
	S = 2;
	#100;


	#100;
	A = 1;
	B = 0;
	S = 2;
	#100;


	#100;
	A = 1;
	B = 1;
	S = 2;
	#100;





	// NOT A TB 
	
	#100;
	A = 0;
	S = 3;
	#100;


	#100;
	A = 1;
	S = 3;
	#100;

*/




	end


endmodule
